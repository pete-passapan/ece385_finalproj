`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/19/2025 11:00:12 AM
// Design Name: 
// Module Name: cottage_cheese
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module cottage_cheese(

    );
    
localparam ADDR_WIDTH = 17; // ceil(log2(76456)) = 17 bits
localparam DEPTH = 76456;

logic [15:0] pcm_rom [DEPTH];



endmodule
