localparam int NUM_LINES = 30;
localparam int NUM_FILTERS = 15;
